module divizor_2(
	input clock, 
	output reg 
); s