module divizor_2(
	input clock, 
	output reg out
); 

always @*
	out = out + 1;

endmodule 